/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`include "mux.v"

`default_nettype none

module tt_um_8_bit_cpu (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire [7:0] a = 8'b01010101;
  wire [7:0] b = 8'b10101010;
  wire [7:0] c = 8'b00001111;
  wire [7:0] d = 8'b11110000;

  wire [1:0] sel = ui_in[1:0];

  wire [7:0] mux_out;

  mux multiplexer (
    .a(a),
    .b(b),
    .c(c),
    .d(d),
    .select(sel),
    .out(mux_out)
  );

  assign uo_out = mux_out;
  assign uio_out = 8'b0;
  assign uio_oe  = 8'b0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, uio_in, 1'b0};

endmodule
